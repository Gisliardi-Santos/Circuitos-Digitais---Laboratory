library IEEE;
use IEEE.std_logic_1164.all;

entity decod_fourSeven is
port(
	a4,a3,a2,a1 : in bit;
	s0,s1,s2,s3,s4,s5,s6 : out bit
	);
end;

architecture main of decod_fourSeven is

begin 
	s0 <= not( a1 ) and not( a3 ) and ( a2 or a4 ) and ( not( a2 ) or not( a4 ) );
	s1 <= not( a1 ) and a2 and ( a3 or a4 ) and ( not( a3 ) or not( a4 ) );
	s2 <= not( a1 ) and not( a2 ) and a3 and not( a4 );
	s3 <= not( a1 ) and (( a2 and a3 and a4 ) or ( a2 and not( a3 ) and not( a4 ) ) or ( not( a2 ) and not( a3 ) and a4 ));
	s4 <= ( not( a1 ) and a4 ) or ( not( a1 ) and a2 and not( a3 ) ) or ( not( a2 ) and not( a3 ) and a4 );
	s5 <= not( a1 ) and ( a3 or a4 ) and ( a3 or not( a4 ) ) and ( not( a2 ) or a4 );
	s6 <= not( a1 ) and (( not( a2 ) and not( a3 ) ) or ( a2 and a3 and a4 ));
end architecture main;